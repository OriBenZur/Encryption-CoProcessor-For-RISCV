// de0cv.v

// Generated using ACDS version 17.0 595

`timescale 1 ps / 1 ps
module de0cv (
		input  wire  clk_clk,       //   clk.clk
		input  wire  reset_reset_n  // reset.reset_n
	);

endmodule
